module SDcardContent(
    input  logic rdclk,
    input  logic [63:0] rdaddr,
    output logic [ 7:0] rddata
);

always @ (posedge rdclk)
    case(rdaddr)
    'h000001B8:rddata=8'h34;
    'h000001B9:rddata=8'h21;
    'h000001BA:rddata=8'h70;
    'h000001BB:rddata=8'h34;
    'h000001BF:rddata=8'h82;
    'h000001C0:rddata=8'h03;
    'h000001C2:rddata=8'h0C;
    'h000001C3:rddata=8'hFE;
    'h000001C4:rddata=8'hFF;
    'h000001C5:rddata=8'hAC;
    'h000001C7:rddata=8'h20;
    'h000001CB:rddata=8'hC0;
    'h000001CC:rddata=8'hE6;
    'h000001FE:rddata=8'h55;
    'h000001FF:rddata=8'hAA;
    'h00400000:rddata=8'hEB;
    'h00400001:rddata=8'h58;
    'h00400002:rddata=8'h90;
    'h00400003:rddata=8'h4D;
    'h00400004:rddata=8'h53;
    'h00400005:rddata=8'h44;
    'h00400006:rddata=8'h4F;
    'h00400007:rddata=8'h53;
    'h00400008:rddata=8'h35;
    'h00400009:rddata=8'h2E;
    'h0040000A:rddata=8'h30;
    'h0040000C:rddata=8'h02;
    'h0040000D:rddata=8'h40;
    'h0040000E:rddata=8'h94;
    'h0040000F:rddata=8'h11;
    'h00400010:rddata=8'h02;
    'h00400015:rddata=8'hF8;
    'h00400018:rddata=8'h3F;
    'h0040001A:rddata=8'hFF;
    'h0040001D:rddata=8'h20;
    'h00400021:rddata=8'hC0;
    'h00400022:rddata=8'hE6;
    'h00400024:rddata=8'h36;
    'h00400025:rddata=8'h07;
    'h0040002C:rddata=8'h02;
    'h00400030:rddata=8'h01;
    'h00400032:rddata=8'h06;
    'h00400040:rddata=8'h80;
    'h00400042:rddata=8'h29;
    'h00400043:rddata=8'h6E;
    'h00400044:rddata=8'hED;
    'h00400045:rddata=8'h87;
    'h00400046:rddata=8'h7E;
    'h00400047:rddata=8'h4E;
    'h00400048:rddata=8'h4F;
    'h00400049:rddata=8'h20;
    'h0040004A:rddata=8'h4E;
    'h0040004B:rddata=8'h41;
    'h0040004C:rddata=8'h4D;
    'h0040004D:rddata=8'h45;
    'h0040004E:rddata=8'h20;
    'h0040004F:rddata=8'h20;
    'h00400050:rddata=8'h20;
    'h00400051:rddata=8'h20;
    'h00400052:rddata=8'h46;
    'h00400053:rddata=8'h41;
    'h00400054:rddata=8'h54;
    'h00400055:rddata=8'h33;
    'h00400056:rddata=8'h32;
    'h00400057:rddata=8'h20;
    'h00400058:rddata=8'h20;
    'h00400059:rddata=8'h20;
    'h0040005A:rddata=8'h33;
    'h0040005B:rddata=8'hC9;
    'h0040005C:rddata=8'h8E;
    'h0040005D:rddata=8'hD1;
    'h0040005E:rddata=8'hBC;
    'h0040005F:rddata=8'hF4;
    'h00400060:rddata=8'h7B;
    'h00400061:rddata=8'h8E;
    'h00400062:rddata=8'hC1;
    'h00400063:rddata=8'h8E;
    'h00400064:rddata=8'hD9;
    'h00400065:rddata=8'hBD;
    'h00400067:rddata=8'h7C;
    'h00400068:rddata=8'h88;
    'h00400069:rddata=8'h56;
    'h0040006A:rddata=8'h40;
    'h0040006B:rddata=8'h88;
    'h0040006C:rddata=8'h4E;
    'h0040006D:rddata=8'h02;
    'h0040006E:rddata=8'h8A;
    'h0040006F:rddata=8'h56;
    'h00400070:rddata=8'h40;
    'h00400071:rddata=8'hB4;
    'h00400072:rddata=8'h41;
    'h00400073:rddata=8'hBB;
    'h00400074:rddata=8'hAA;
    'h00400075:rddata=8'h55;
    'h00400076:rddata=8'hCD;
    'h00400077:rddata=8'h13;
    'h00400078:rddata=8'h72;
    'h00400079:rddata=8'h10;
    'h0040007A:rddata=8'h81;
    'h0040007B:rddata=8'hFB;
    'h0040007C:rddata=8'h55;
    'h0040007D:rddata=8'hAA;
    'h0040007E:rddata=8'h75;
    'h0040007F:rddata=8'h0A;
    'h00400080:rddata=8'hF6;
    'h00400081:rddata=8'hC1;
    'h00400082:rddata=8'h01;
    'h00400083:rddata=8'h74;
    'h00400084:rddata=8'h05;
    'h00400085:rddata=8'hFE;
    'h00400086:rddata=8'h46;
    'h00400087:rddata=8'h02;
    'h00400088:rddata=8'hEB;
    'h00400089:rddata=8'h2D;
    'h0040008A:rddata=8'h8A;
    'h0040008B:rddata=8'h56;
    'h0040008C:rddata=8'h40;
    'h0040008D:rddata=8'hB4;
    'h0040008E:rddata=8'h08;
    'h0040008F:rddata=8'hCD;
    'h00400090:rddata=8'h13;
    'h00400091:rddata=8'h73;
    'h00400092:rddata=8'h05;
    'h00400093:rddata=8'hB9;
    'h00400094:rddata=8'hFF;
    'h00400095:rddata=8'hFF;
    'h00400096:rddata=8'h8A;
    'h00400097:rddata=8'hF1;
    'h00400098:rddata=8'h66;
    'h00400099:rddata=8'h0F;
    'h0040009A:rddata=8'hB6;
    'h0040009B:rddata=8'hC6;
    'h0040009C:rddata=8'h40;
    'h0040009D:rddata=8'h66;
    'h0040009E:rddata=8'h0F;
    'h0040009F:rddata=8'hB6;
    'h004000A0:rddata=8'hD1;
    'h004000A1:rddata=8'h80;
    'h004000A2:rddata=8'hE2;
    'h004000A3:rddata=8'h3F;
    'h004000A4:rddata=8'hF7;
    'h004000A5:rddata=8'hE2;
    'h004000A6:rddata=8'h86;
    'h004000A7:rddata=8'hCD;
    'h004000A8:rddata=8'hC0;
    'h004000A9:rddata=8'hED;
    'h004000AA:rddata=8'h06;
    'h004000AB:rddata=8'h41;
    'h004000AC:rddata=8'h66;
    'h004000AD:rddata=8'h0F;
    'h004000AE:rddata=8'hB7;
    'h004000AF:rddata=8'hC9;
    'h004000B0:rddata=8'h66;
    'h004000B1:rddata=8'hF7;
    'h004000B2:rddata=8'hE1;
    'h004000B3:rddata=8'h66;
    'h004000B4:rddata=8'h89;
    'h004000B5:rddata=8'h46;
    'h004000B6:rddata=8'hF8;
    'h004000B7:rddata=8'h83;
    'h004000B8:rddata=8'h7E;
    'h004000B9:rddata=8'h16;
    'h004000BB:rddata=8'h75;
    'h004000BC:rddata=8'h39;
    'h004000BD:rddata=8'h83;
    'h004000BE:rddata=8'h7E;
    'h004000BF:rddata=8'h2A;
    'h004000C1:rddata=8'h77;
    'h004000C2:rddata=8'h33;
    'h004000C3:rddata=8'h66;
    'h004000C4:rddata=8'h8B;
    'h004000C5:rddata=8'h46;
    'h004000C6:rddata=8'h1C;
    'h004000C7:rddata=8'h66;
    'h004000C8:rddata=8'h83;
    'h004000C9:rddata=8'hC0;
    'h004000CA:rddata=8'h0C;
    'h004000CB:rddata=8'hBB;
    'h004000CD:rddata=8'h80;
    'h004000CE:rddata=8'hB9;
    'h004000CF:rddata=8'h01;
    'h004000D1:rddata=8'hE8;
    'h004000D2:rddata=8'h2C;
    'h004000D4:rddata=8'hE9;
    'h004000D5:rddata=8'hA8;
    'h004000D6:rddata=8'h03;
    'h004000D7:rddata=8'hA1;
    'h004000D8:rddata=8'hF8;
    'h004000D9:rddata=8'h7D;
    'h004000DA:rddata=8'h80;
    'h004000DB:rddata=8'hC4;
    'h004000DC:rddata=8'h7C;
    'h004000DD:rddata=8'h8B;
    'h004000DE:rddata=8'hF0;
    'h004000DF:rddata=8'hAC;
    'h004000E0:rddata=8'h84;
    'h004000E1:rddata=8'hC0;
    'h004000E2:rddata=8'h74;
    'h004000E3:rddata=8'h17;
    'h004000E4:rddata=8'h3C;
    'h004000E5:rddata=8'hFF;
    'h004000E6:rddata=8'h74;
    'h004000E7:rddata=8'h09;
    'h004000E8:rddata=8'hB4;
    'h004000E9:rddata=8'h0E;
    'h004000EA:rddata=8'hBB;
    'h004000EB:rddata=8'h07;
    'h004000ED:rddata=8'hCD;
    'h004000EE:rddata=8'h10;
    'h004000EF:rddata=8'hEB;
    'h004000F0:rddata=8'hEE;
    'h004000F1:rddata=8'hA1;
    'h004000F2:rddata=8'hFA;
    'h004000F3:rddata=8'h7D;
    'h004000F4:rddata=8'hEB;
    'h004000F5:rddata=8'hE4;
    'h004000F6:rddata=8'hA1;
    'h004000F7:rddata=8'h7D;
    'h004000F8:rddata=8'h80;
    'h004000F9:rddata=8'hEB;
    'h004000FA:rddata=8'hDF;
    'h004000FB:rddata=8'h98;
    'h004000FC:rddata=8'hCD;
    'h004000FD:rddata=8'h16;
    'h004000FE:rddata=8'hCD;
    'h004000FF:rddata=8'h19;
    'h00400100:rddata=8'h66;
    'h00400101:rddata=8'h60;
    'h00400102:rddata=8'h80;
    'h00400103:rddata=8'h7E;
    'h00400104:rddata=8'h02;
    'h00400106:rddata=8'h0F;
    'h00400107:rddata=8'h84;
    'h00400108:rddata=8'h20;
    'h0040010A:rddata=8'h66;
    'h0040010B:rddata=8'h6A;
    'h0040010D:rddata=8'h66;
    'h0040010E:rddata=8'h50;
    'h0040010F:rddata=8'h06;
    'h00400110:rddata=8'h53;
    'h00400111:rddata=8'h66;
    'h00400112:rddata=8'h68;
    'h00400113:rddata=8'h10;
    'h00400115:rddata=8'h01;
    'h00400117:rddata=8'hB4;
    'h00400118:rddata=8'h42;
    'h00400119:rddata=8'h8A;
    'h0040011A:rddata=8'h56;
    'h0040011B:rddata=8'h40;
    'h0040011C:rddata=8'h8B;
    'h0040011D:rddata=8'hF4;
    'h0040011E:rddata=8'hCD;
    'h0040011F:rddata=8'h13;
    'h00400120:rddata=8'h66;
    'h00400121:rddata=8'h58;
    'h00400122:rddata=8'h66;
    'h00400123:rddata=8'h58;
    'h00400124:rddata=8'h66;
    'h00400125:rddata=8'h58;
    'h00400126:rddata=8'h66;
    'h00400127:rddata=8'h58;
    'h00400128:rddata=8'hEB;
    'h00400129:rddata=8'h33;
    'h0040012A:rddata=8'h66;
    'h0040012B:rddata=8'h3B;
    'h0040012C:rddata=8'h46;
    'h0040012D:rddata=8'hF8;
    'h0040012E:rddata=8'h72;
    'h0040012F:rddata=8'h03;
    'h00400130:rddata=8'hF9;
    'h00400131:rddata=8'hEB;
    'h00400132:rddata=8'h2A;
    'h00400133:rddata=8'h66;
    'h00400134:rddata=8'h33;
    'h00400135:rddata=8'hD2;
    'h00400136:rddata=8'h66;
    'h00400137:rddata=8'h0F;
    'h00400138:rddata=8'hB7;
    'h00400139:rddata=8'h4E;
    'h0040013A:rddata=8'h18;
    'h0040013B:rddata=8'h66;
    'h0040013C:rddata=8'hF7;
    'h0040013D:rddata=8'hF1;
    'h0040013E:rddata=8'hFE;
    'h0040013F:rddata=8'hC2;
    'h00400140:rddata=8'h8A;
    'h00400141:rddata=8'hCA;
    'h00400142:rddata=8'h66;
    'h00400143:rddata=8'h8B;
    'h00400144:rddata=8'hD0;
    'h00400145:rddata=8'h66;
    'h00400146:rddata=8'hC1;
    'h00400147:rddata=8'hEA;
    'h00400148:rddata=8'h10;
    'h00400149:rddata=8'hF7;
    'h0040014A:rddata=8'h76;
    'h0040014B:rddata=8'h1A;
    'h0040014C:rddata=8'h86;
    'h0040014D:rddata=8'hD6;
    'h0040014E:rddata=8'h8A;
    'h0040014F:rddata=8'h56;
    'h00400150:rddata=8'h40;
    'h00400151:rddata=8'h8A;
    'h00400152:rddata=8'hE8;
    'h00400153:rddata=8'hC0;
    'h00400154:rddata=8'hE4;
    'h00400155:rddata=8'h06;
    'h00400156:rddata=8'h0A;
    'h00400157:rddata=8'hCC;
    'h00400158:rddata=8'hB8;
    'h00400159:rddata=8'h01;
    'h0040015A:rddata=8'h02;
    'h0040015B:rddata=8'hCD;
    'h0040015C:rddata=8'h13;
    'h0040015D:rddata=8'h66;
    'h0040015E:rddata=8'h61;
    'h0040015F:rddata=8'h0F;
    'h00400160:rddata=8'h82;
    'h00400161:rddata=8'h74;
    'h00400162:rddata=8'hFF;
    'h00400163:rddata=8'h81;
    'h00400164:rddata=8'hC3;
    'h00400166:rddata=8'h02;
    'h00400167:rddata=8'h66;
    'h00400168:rddata=8'h40;
    'h00400169:rddata=8'h49;
    'h0040016A:rddata=8'h75;
    'h0040016B:rddata=8'h94;
    'h0040016C:rddata=8'hC3;
    'h0040016D:rddata=8'h42;
    'h0040016E:rddata=8'h4F;
    'h0040016F:rddata=8'h4F;
    'h00400170:rddata=8'h54;
    'h00400171:rddata=8'h4D;
    'h00400172:rddata=8'h47;
    'h00400173:rddata=8'h52;
    'h00400174:rddata=8'h20;
    'h00400175:rddata=8'h20;
    'h00400176:rddata=8'h20;
    'h00400177:rddata=8'h20;
    'h004001AC:rddata=8'h0D;
    'h004001AD:rddata=8'h0A;
    'h004001AE:rddata=8'h44;
    'h004001AF:rddata=8'h69;
    'h004001B0:rddata=8'h73;
    'h004001B1:rddata=8'h6B;
    'h004001B2:rddata=8'h20;
    'h004001B3:rddata=8'h65;
    'h004001B4:rddata=8'h72;
    'h004001B5:rddata=8'h72;
    'h004001B6:rddata=8'h6F;
    'h004001B7:rddata=8'h72;
    'h004001B8:rddata=8'hFF;
    'h004001B9:rddata=8'h0D;
    'h004001BA:rddata=8'h0A;
    'h004001BB:rddata=8'h50;
    'h004001BC:rddata=8'h72;
    'h004001BD:rddata=8'h65;
    'h004001BE:rddata=8'h73;
    'h004001BF:rddata=8'h73;
    'h004001C0:rddata=8'h20;
    'h004001C1:rddata=8'h61;
    'h004001C2:rddata=8'h6E;
    'h004001C3:rddata=8'h79;
    'h004001C4:rddata=8'h20;
    'h004001C5:rddata=8'h6B;
    'h004001C6:rddata=8'h65;
    'h004001C7:rddata=8'h79;
    'h004001C8:rddata=8'h20;
    'h004001C9:rddata=8'h74;
    'h004001CA:rddata=8'h6F;
    'h004001CB:rddata=8'h20;
    'h004001CC:rddata=8'h72;
    'h004001CD:rddata=8'h65;
    'h004001CE:rddata=8'h73;
    'h004001CF:rddata=8'h74;
    'h004001D0:rddata=8'h61;
    'h004001D1:rddata=8'h72;
    'h004001D2:rddata=8'h74;
    'h004001D3:rddata=8'h0D;
    'h004001D4:rddata=8'h0A;
    'h004001F8:rddata=8'hAC;
    'h004001F9:rddata=8'h01;
    'h004001FA:rddata=8'hB9;
    'h004001FB:rddata=8'h01;
    'h004001FE:rddata=8'h55;
    'h004001FF:rddata=8'hAA;
    'h00400200:rddata=8'h52;
    'h00400201:rddata=8'h52;
    'h00400202:rddata=8'h61;
    'h00400203:rddata=8'h41;
    'h004003E4:rddata=8'h72;
    'h004003E5:rddata=8'h72;
    'h004003E6:rddata=8'h41;
    'h004003E7:rddata=8'h61;
    'h004003E8:rddata=8'h7B;
    'h004003E9:rddata=8'h9A;
    'h004003EA:rddata=8'h03;
    'h004003EC:rddata=8'h07;
    'h004003FE:rddata=8'h55;
    'h004003FF:rddata=8'hAA;
    'h004005FE:rddata=8'h55;
    'h004005FF:rddata=8'hAA;
    'h00400C00:rddata=8'hEB;
    'h00400C01:rddata=8'h58;
    'h00400C02:rddata=8'h90;
    'h00400C03:rddata=8'h4D;
    'h00400C04:rddata=8'h53;
    'h00400C05:rddata=8'h44;
    'h00400C06:rddata=8'h4F;
    'h00400C07:rddata=8'h53;
    'h00400C08:rddata=8'h35;
    'h00400C09:rddata=8'h2E;
    'h00400C0A:rddata=8'h30;
    'h00400C0C:rddata=8'h02;
    'h00400C0D:rddata=8'h40;
    'h00400C0E:rddata=8'h94;
    'h00400C0F:rddata=8'h11;
    'h00400C10:rddata=8'h02;
    'h00400C15:rddata=8'hF8;
    'h00400C18:rddata=8'h3F;
    'h00400C1A:rddata=8'hFF;
    'h00400C1D:rddata=8'h20;
    'h00400C21:rddata=8'hC0;
    'h00400C22:rddata=8'hE6;
    'h00400C24:rddata=8'h36;
    'h00400C25:rddata=8'h07;
    'h00400C2C:rddata=8'h02;
    'h00400C30:rddata=8'h01;
    'h00400C32:rddata=8'h06;
    'h00400C40:rddata=8'h80;
    'h00400C42:rddata=8'h29;
    'h00400C43:rddata=8'h6E;
    'h00400C44:rddata=8'hED;
    'h00400C45:rddata=8'h87;
    'h00400C46:rddata=8'h7E;
    'h00400C47:rddata=8'h4E;
    'h00400C48:rddata=8'h4F;
    'h00400C49:rddata=8'h20;
    'h00400C4A:rddata=8'h4E;
    'h00400C4B:rddata=8'h41;
    'h00400C4C:rddata=8'h4D;
    'h00400C4D:rddata=8'h45;
    'h00400C4E:rddata=8'h20;
    'h00400C4F:rddata=8'h20;
    'h00400C50:rddata=8'h20;
    'h00400C51:rddata=8'h20;
    'h00400C52:rddata=8'h46;
    'h00400C53:rddata=8'h41;
    'h00400C54:rddata=8'h54;
    'h00400C55:rddata=8'h33;
    'h00400C56:rddata=8'h32;
    'h00400C57:rddata=8'h20;
    'h00400C58:rddata=8'h20;
    'h00400C59:rddata=8'h20;
    'h00400C5A:rddata=8'h33;
    'h00400C5B:rddata=8'hC9;
    'h00400C5C:rddata=8'h8E;
    'h00400C5D:rddata=8'hD1;
    'h00400C5E:rddata=8'hBC;
    'h00400C5F:rddata=8'hF4;
    'h00400C60:rddata=8'h7B;
    'h00400C61:rddata=8'h8E;
    'h00400C62:rddata=8'hC1;
    'h00400C63:rddata=8'h8E;
    'h00400C64:rddata=8'hD9;
    'h00400C65:rddata=8'hBD;
    'h00400C67:rddata=8'h7C;
    'h00400C68:rddata=8'h88;
    'h00400C69:rddata=8'h56;
    'h00400C6A:rddata=8'h40;
    'h00400C6B:rddata=8'h88;
    'h00400C6C:rddata=8'h4E;
    'h00400C6D:rddata=8'h02;
    'h00400C6E:rddata=8'h8A;
    'h00400C6F:rddata=8'h56;
    'h00400C70:rddata=8'h40;
    'h00400C71:rddata=8'hB4;
    'h00400C72:rddata=8'h41;
    'h00400C73:rddata=8'hBB;
    'h00400C74:rddata=8'hAA;
    'h00400C75:rddata=8'h55;
    'h00400C76:rddata=8'hCD;
    'h00400C77:rddata=8'h13;
    'h00400C78:rddata=8'h72;
    'h00400C79:rddata=8'h10;
    'h00400C7A:rddata=8'h81;
    'h00400C7B:rddata=8'hFB;
    'h00400C7C:rddata=8'h55;
    'h00400C7D:rddata=8'hAA;
    'h00400C7E:rddata=8'h75;
    'h00400C7F:rddata=8'h0A;
    'h00400C80:rddata=8'hF6;
    'h00400C81:rddata=8'hC1;
    'h00400C82:rddata=8'h01;
    'h00400C83:rddata=8'h74;
    'h00400C84:rddata=8'h05;
    'h00400C85:rddata=8'hFE;
    'h00400C86:rddata=8'h46;
    'h00400C87:rddata=8'h02;
    'h00400C88:rddata=8'hEB;
    'h00400C89:rddata=8'h2D;
    'h00400C8A:rddata=8'h8A;
    'h00400C8B:rddata=8'h56;
    'h00400C8C:rddata=8'h40;
    'h00400C8D:rddata=8'hB4;
    'h00400C8E:rddata=8'h08;
    'h00400C8F:rddata=8'hCD;
    'h00400C90:rddata=8'h13;
    'h00400C91:rddata=8'h73;
    'h00400C92:rddata=8'h05;
    'h00400C93:rddata=8'hB9;
    'h00400C94:rddata=8'hFF;
    'h00400C95:rddata=8'hFF;
    'h00400C96:rddata=8'h8A;
    'h00400C97:rddata=8'hF1;
    'h00400C98:rddata=8'h66;
    'h00400C99:rddata=8'h0F;
    'h00400C9A:rddata=8'hB6;
    'h00400C9B:rddata=8'hC6;
    'h00400C9C:rddata=8'h40;
    'h00400C9D:rddata=8'h66;
    'h00400C9E:rddata=8'h0F;
    'h00400C9F:rddata=8'hB6;
    'h00400CA0:rddata=8'hD1;
    'h00400CA1:rddata=8'h80;
    'h00400CA2:rddata=8'hE2;
    'h00400CA3:rddata=8'h3F;
    'h00400CA4:rddata=8'hF7;
    'h00400CA5:rddata=8'hE2;
    'h00400CA6:rddata=8'h86;
    'h00400CA7:rddata=8'hCD;
    'h00400CA8:rddata=8'hC0;
    'h00400CA9:rddata=8'hED;
    'h00400CAA:rddata=8'h06;
    'h00400CAB:rddata=8'h41;
    'h00400CAC:rddata=8'h66;
    'h00400CAD:rddata=8'h0F;
    'h00400CAE:rddata=8'hB7;
    'h00400CAF:rddata=8'hC9;
    'h00400CB0:rddata=8'h66;
    'h00400CB1:rddata=8'hF7;
    'h00400CB2:rddata=8'hE1;
    'h00400CB3:rddata=8'h66;
    'h00400CB4:rddata=8'h89;
    'h00400CB5:rddata=8'h46;
    'h00400CB6:rddata=8'hF8;
    'h00400CB7:rddata=8'h83;
    'h00400CB8:rddata=8'h7E;
    'h00400CB9:rddata=8'h16;
    'h00400CBB:rddata=8'h75;
    'h00400CBC:rddata=8'h39;
    'h00400CBD:rddata=8'h83;
    'h00400CBE:rddata=8'h7E;
    'h00400CBF:rddata=8'h2A;
    'h00400CC1:rddata=8'h77;
    'h00400CC2:rddata=8'h33;
    'h00400CC3:rddata=8'h66;
    'h00400CC4:rddata=8'h8B;
    'h00400CC5:rddata=8'h46;
    'h00400CC6:rddata=8'h1C;
    'h00400CC7:rddata=8'h66;
    'h00400CC8:rddata=8'h83;
    'h00400CC9:rddata=8'hC0;
    'h00400CCA:rddata=8'h0C;
    'h00400CCB:rddata=8'hBB;
    'h00400CCD:rddata=8'h80;
    'h00400CCE:rddata=8'hB9;
    'h00400CCF:rddata=8'h01;
    'h00400CD1:rddata=8'hE8;
    'h00400CD2:rddata=8'h2C;
    'h00400CD4:rddata=8'hE9;
    'h00400CD5:rddata=8'hA8;
    'h00400CD6:rddata=8'h03;
    'h00400CD7:rddata=8'hA1;
    'h00400CD8:rddata=8'hF8;
    'h00400CD9:rddata=8'h7D;
    'h00400CDA:rddata=8'h80;
    'h00400CDB:rddata=8'hC4;
    'h00400CDC:rddata=8'h7C;
    'h00400CDD:rddata=8'h8B;
    'h00400CDE:rddata=8'hF0;
    'h00400CDF:rddata=8'hAC;
    'h00400CE0:rddata=8'h84;
    'h00400CE1:rddata=8'hC0;
    'h00400CE2:rddata=8'h74;
    'h00400CE3:rddata=8'h17;
    'h00400CE4:rddata=8'h3C;
    'h00400CE5:rddata=8'hFF;
    'h00400CE6:rddata=8'h74;
    'h00400CE7:rddata=8'h09;
    'h00400CE8:rddata=8'hB4;
    'h00400CE9:rddata=8'h0E;
    'h00400CEA:rddata=8'hBB;
    'h00400CEB:rddata=8'h07;
    'h00400CED:rddata=8'hCD;
    'h00400CEE:rddata=8'h10;
    'h00400CEF:rddata=8'hEB;
    'h00400CF0:rddata=8'hEE;
    'h00400CF1:rddata=8'hA1;
    'h00400CF2:rddata=8'hFA;
    'h00400CF3:rddata=8'h7D;
    'h00400CF4:rddata=8'hEB;
    'h00400CF5:rddata=8'hE4;
    'h00400CF6:rddata=8'hA1;
    'h00400CF7:rddata=8'h7D;
    'h00400CF8:rddata=8'h80;
    'h00400CF9:rddata=8'hEB;
    'h00400CFA:rddata=8'hDF;
    'h00400CFB:rddata=8'h98;
    'h00400CFC:rddata=8'hCD;
    'h00400CFD:rddata=8'h16;
    'h00400CFE:rddata=8'hCD;
    'h00400CFF:rddata=8'h19;
    'h00400D00:rddata=8'h66;
    'h00400D01:rddata=8'h60;
    'h00400D02:rddata=8'h80;
    'h00400D03:rddata=8'h7E;
    'h00400D04:rddata=8'h02;
    'h00400D06:rddata=8'h0F;
    'h00400D07:rddata=8'h84;
    'h00400D08:rddata=8'h20;
    'h00400D0A:rddata=8'h66;
    'h00400D0B:rddata=8'h6A;
    'h00400D0D:rddata=8'h66;
    'h00400D0E:rddata=8'h50;
    'h00400D0F:rddata=8'h06;
    'h00400D10:rddata=8'h53;
    'h00400D11:rddata=8'h66;
    'h00400D12:rddata=8'h68;
    'h00400D13:rddata=8'h10;
    'h00400D15:rddata=8'h01;
    'h00400D17:rddata=8'hB4;
    'h00400D18:rddata=8'h42;
    'h00400D19:rddata=8'h8A;
    'h00400D1A:rddata=8'h56;
    'h00400D1B:rddata=8'h40;
    'h00400D1C:rddata=8'h8B;
    'h00400D1D:rddata=8'hF4;
    'h00400D1E:rddata=8'hCD;
    'h00400D1F:rddata=8'h13;
    'h00400D20:rddata=8'h66;
    'h00400D21:rddata=8'h58;
    'h00400D22:rddata=8'h66;
    'h00400D23:rddata=8'h58;
    'h00400D24:rddata=8'h66;
    'h00400D25:rddata=8'h58;
    'h00400D26:rddata=8'h66;
    'h00400D27:rddata=8'h58;
    'h00400D28:rddata=8'hEB;
    'h00400D29:rddata=8'h33;
    'h00400D2A:rddata=8'h66;
    'h00400D2B:rddata=8'h3B;
    'h00400D2C:rddata=8'h46;
    'h00400D2D:rddata=8'hF8;
    'h00400D2E:rddata=8'h72;
    'h00400D2F:rddata=8'h03;
    'h00400D30:rddata=8'hF9;
    'h00400D31:rddata=8'hEB;
    'h00400D32:rddata=8'h2A;
    'h00400D33:rddata=8'h66;
    'h00400D34:rddata=8'h33;
    'h00400D35:rddata=8'hD2;
    'h00400D36:rddata=8'h66;
    'h00400D37:rddata=8'h0F;
    'h00400D38:rddata=8'hB7;
    'h00400D39:rddata=8'h4E;
    'h00400D3A:rddata=8'h18;
    'h00400D3B:rddata=8'h66;
    'h00400D3C:rddata=8'hF7;
    'h00400D3D:rddata=8'hF1;
    'h00400D3E:rddata=8'hFE;
    'h00400D3F:rddata=8'hC2;
    'h00400D40:rddata=8'h8A;
    'h00400D41:rddata=8'hCA;
    'h00400D42:rddata=8'h66;
    'h00400D43:rddata=8'h8B;
    'h00400D44:rddata=8'hD0;
    'h00400D45:rddata=8'h66;
    'h00400D46:rddata=8'hC1;
    'h00400D47:rddata=8'hEA;
    'h00400D48:rddata=8'h10;
    'h00400D49:rddata=8'hF7;
    'h00400D4A:rddata=8'h76;
    'h00400D4B:rddata=8'h1A;
    'h00400D4C:rddata=8'h86;
    'h00400D4D:rddata=8'hD6;
    'h00400D4E:rddata=8'h8A;
    'h00400D4F:rddata=8'h56;
    'h00400D50:rddata=8'h40;
    'h00400D51:rddata=8'h8A;
    'h00400D52:rddata=8'hE8;
    'h00400D53:rddata=8'hC0;
    'h00400D54:rddata=8'hE4;
    'h00400D55:rddata=8'h06;
    'h00400D56:rddata=8'h0A;
    'h00400D57:rddata=8'hCC;
    'h00400D58:rddata=8'hB8;
    'h00400D59:rddata=8'h01;
    'h00400D5A:rddata=8'h02;
    'h00400D5B:rddata=8'hCD;
    'h00400D5C:rddata=8'h13;
    'h00400D5D:rddata=8'h66;
    'h00400D5E:rddata=8'h61;
    'h00400D5F:rddata=8'h0F;
    'h00400D60:rddata=8'h82;
    'h00400D61:rddata=8'h74;
    'h00400D62:rddata=8'hFF;
    'h00400D63:rddata=8'h81;
    'h00400D64:rddata=8'hC3;
    'h00400D66:rddata=8'h02;
    'h00400D67:rddata=8'h66;
    'h00400D68:rddata=8'h40;
    'h00400D69:rddata=8'h49;
    'h00400D6A:rddata=8'h75;
    'h00400D6B:rddata=8'h94;
    'h00400D6C:rddata=8'hC3;
    'h00400D6D:rddata=8'h42;
    'h00400D6E:rddata=8'h4F;
    'h00400D6F:rddata=8'h4F;
    'h00400D70:rddata=8'h54;
    'h00400D71:rddata=8'h4D;
    'h00400D72:rddata=8'h47;
    'h00400D73:rddata=8'h52;
    'h00400D74:rddata=8'h20;
    'h00400D75:rddata=8'h20;
    'h00400D76:rddata=8'h20;
    'h00400D77:rddata=8'h20;
    'h00400DAC:rddata=8'h0D;
    'h00400DAD:rddata=8'h0A;
    'h00400DAE:rddata=8'h44;
    'h00400DAF:rddata=8'h69;
    'h00400DB0:rddata=8'h73;
    'h00400DB1:rddata=8'h6B;
    'h00400DB2:rddata=8'h20;
    'h00400DB3:rddata=8'h65;
    'h00400DB4:rddata=8'h72;
    'h00400DB5:rddata=8'h72;
    'h00400DB6:rddata=8'h6F;
    'h00400DB7:rddata=8'h72;
    'h00400DB8:rddata=8'hFF;
    'h00400DB9:rddata=8'h0D;
    'h00400DBA:rddata=8'h0A;
    'h00400DBB:rddata=8'h50;
    'h00400DBC:rddata=8'h72;
    'h00400DBD:rddata=8'h65;
    'h00400DBE:rddata=8'h73;
    'h00400DBF:rddata=8'h73;
    'h00400DC0:rddata=8'h20;
    'h00400DC1:rddata=8'h61;
    'h00400DC2:rddata=8'h6E;
    'h00400DC3:rddata=8'h79;
    'h00400DC4:rddata=8'h20;
    'h00400DC5:rddata=8'h6B;
    'h00400DC6:rddata=8'h65;
    'h00400DC7:rddata=8'h79;
    'h00400DC8:rddata=8'h20;
    'h00400DC9:rddata=8'h74;
    'h00400DCA:rddata=8'h6F;
    'h00400DCB:rddata=8'h20;
    'h00400DCC:rddata=8'h72;
    'h00400DCD:rddata=8'h65;
    'h00400DCE:rddata=8'h73;
    'h00400DCF:rddata=8'h74;
    'h00400DD0:rddata=8'h61;
    'h00400DD1:rddata=8'h72;
    'h00400DD2:rddata=8'h74;
    'h00400DD3:rddata=8'h0D;
    'h00400DD4:rddata=8'h0A;
    'h00400DF8:rddata=8'hAC;
    'h00400DF9:rddata=8'h01;
    'h00400DFA:rddata=8'hB9;
    'h00400DFB:rddata=8'h01;
    'h00400DFE:rddata=8'h55;
    'h00400DFF:rddata=8'hAA;
    'h00400E00:rddata=8'h52;
    'h00400E01:rddata=8'h52;
    'h00400E02:rddata=8'h61;
    'h00400E03:rddata=8'h41;
    'h00400FE4:rddata=8'h72;
    'h00400FE5:rddata=8'h72;
    'h00400FE6:rddata=8'h41;
    'h00400FE7:rddata=8'h61;
    'h00400FE8:rddata=8'hFF;
    'h00400FE9:rddata=8'hFF;
    'h00400FEA:rddata=8'hFF;
    'h00400FEB:rddata=8'hFF;
    'h00400FEC:rddata=8'h02;
    'h00400FFE:rddata=8'h55;
    'h00400FFF:rddata=8'hAA;
    'h004011FE:rddata=8'h55;
    'h004011FF:rddata=8'hAA;
    'h00401800:rddata=8'h0D;
    'h00401801:rddata=8'h0A;
    'h00401802:rddata=8'h41;
    'h00401803:rddata=8'h6E;
    'h00401804:rddata=8'h20;
    'h00401805:rddata=8'h6F;
    'h00401806:rddata=8'h70;
    'h00401807:rddata=8'h65;
    'h00401808:rddata=8'h72;
    'h00401809:rddata=8'h61;
    'h0040180A:rddata=8'h74;
    'h0040180B:rddata=8'h69;
    'h0040180C:rddata=8'h6E;
    'h0040180D:rddata=8'h67;
    'h0040180E:rddata=8'h20;
    'h0040180F:rddata=8'h73;
    'h00401810:rddata=8'h79;
    'h00401811:rddata=8'h73;
    'h00401812:rddata=8'h74;
    'h00401813:rddata=8'h65;
    'h00401814:rddata=8'h6D;
    'h00401815:rddata=8'h20;
    'h00401816:rddata=8'h77;
    'h00401817:rddata=8'h61;
    'h00401818:rddata=8'h73;
    'h00401819:rddata=8'h6E;
    'h0040181A:rddata=8'h27;
    'h0040181B:rddata=8'h74;
    'h0040181C:rddata=8'h20;
    'h0040181D:rddata=8'h66;
    'h0040181E:rddata=8'h6F;
    'h0040181F:rddata=8'h75;
    'h00401820:rddata=8'h6E;
    'h00401821:rddata=8'h64;
    'h00401822:rddata=8'h2E;
    'h00401823:rddata=8'h20;
    'h00401824:rddata=8'h54;
    'h00401825:rddata=8'h72;
    'h00401826:rddata=8'h79;
    'h00401827:rddata=8'h20;
    'h00401828:rddata=8'h64;
    'h00401829:rddata=8'h69;
    'h0040182A:rddata=8'h73;
    'h0040182B:rddata=8'h63;
    'h0040182C:rddata=8'h6F;
    'h0040182D:rddata=8'h6E;
    'h0040182E:rddata=8'h6E;
    'h0040182F:rddata=8'h65;
    'h00401830:rddata=8'h63;
    'h00401831:rddata=8'h74;
    'h00401832:rddata=8'h69;
    'h00401833:rddata=8'h6E;
    'h00401834:rddata=8'h67;
    'h00401835:rddata=8'h20;
    'h00401836:rddata=8'h61;
    'h00401837:rddata=8'h6E;
    'h00401838:rddata=8'h79;
    'h00401839:rddata=8'h20;
    'h0040183A:rddata=8'h64;
    'h0040183B:rddata=8'h72;
    'h0040183C:rddata=8'h69;
    'h0040183D:rddata=8'h76;
    'h0040183E:rddata=8'h65;
    'h0040183F:rddata=8'h73;
    'h00401840:rddata=8'h20;
    'h00401841:rddata=8'h74;
    'h00401842:rddata=8'h68;
    'h00401843:rddata=8'h61;
    'h00401844:rddata=8'h74;
    'h00401845:rddata=8'h20;
    'h00401846:rddata=8'h64;
    'h00401847:rddata=8'h6F;
    'h00401848:rddata=8'h6E;
    'h00401849:rddata=8'h27;
    'h0040184A:rddata=8'h74;
    'h0040184B:rddata=8'h0D;
    'h0040184C:rddata=8'h0A;
    'h0040184D:rddata=8'h63;
    'h0040184E:rddata=8'h6F;
    'h0040184F:rddata=8'h6E;
    'h00401850:rddata=8'h74;
    'h00401851:rddata=8'h61;
    'h00401852:rddata=8'h69;
    'h00401853:rddata=8'h6E;
    'h00401854:rddata=8'h20;
    'h00401855:rddata=8'h61;
    'h00401856:rddata=8'h6E;
    'h00401857:rddata=8'h20;
    'h00401858:rddata=8'h6F;
    'h00401859:rddata=8'h70;
    'h0040185A:rddata=8'h65;
    'h0040185B:rddata=8'h72;
    'h0040185C:rddata=8'h61;
    'h0040185D:rddata=8'h74;
    'h0040185E:rddata=8'h69;
    'h0040185F:rddata=8'h6E;
    'h00401860:rddata=8'h67;
    'h00401861:rddata=8'h20;
    'h00401862:rddata=8'h73;
    'h00401863:rddata=8'h79;
    'h00401864:rddata=8'h73;
    'h00401865:rddata=8'h74;
    'h00401866:rddata=8'h65;
    'h00401867:rddata=8'h6D;
    'h00401868:rddata=8'h2E;
    'h00401869:rddata=8'hFF;
    'h0040187E:rddata=8'h04;
    'h0040187F:rddata=8'h66;
    'h00401880:rddata=8'h0F;
    'h00401881:rddata=8'hB6;
    'h00401882:rddata=8'h46;
    'h00401883:rddata=8'h10;
    'h00401884:rddata=8'h66;
    'h00401885:rddata=8'h8B;
    'h00401886:rddata=8'h4E;
    'h00401887:rddata=8'h24;
    'h00401888:rddata=8'h66;
    'h00401889:rddata=8'hF7;
    'h0040188A:rddata=8'hE1;
    'h0040188B:rddata=8'h66;
    'h0040188C:rddata=8'h03;
    'h0040188D:rddata=8'h46;
    'h0040188E:rddata=8'h1C;
    'h0040188F:rddata=8'h66;
    'h00401890:rddata=8'h0F;
    'h00401891:rddata=8'hB7;
    'h00401892:rddata=8'h56;
    'h00401893:rddata=8'h0E;
    'h00401894:rddata=8'h66;
    'h00401895:rddata=8'h03;
    'h00401896:rddata=8'hC2;
    'h00401897:rddata=8'h66;
    'h00401898:rddata=8'h89;
    'h00401899:rddata=8'h46;
    'h0040189A:rddata=8'hFC;
    'h0040189B:rddata=8'h66;
    'h0040189C:rddata=8'hC7;
    'h0040189D:rddata=8'h46;
    'h0040189E:rddata=8'hF4;
    'h0040189F:rddata=8'hFF;
    'h004018A0:rddata=8'hFF;
    'h004018A1:rddata=8'hFF;
    'h004018A2:rddata=8'hFF;
    'h004018A3:rddata=8'h66;
    'h004018A4:rddata=8'h8B;
    'h004018A5:rddata=8'h46;
    'h004018A6:rddata=8'h2C;
    'h004018A7:rddata=8'h66;
    'h004018A8:rddata=8'h83;
    'h004018A9:rddata=8'hF8;
    'h004018AA:rddata=8'h02;
    'h004018AB:rddata=8'h0F;
    'h004018AC:rddata=8'h82;
    'h004018AD:rddata=8'h47;
    'h004018AE:rddata=8'hFC;
    'h004018AF:rddata=8'h66;
    'h004018B0:rddata=8'h3D;
    'h004018B1:rddata=8'hF8;
    'h004018B2:rddata=8'hFF;
    'h004018B3:rddata=8'hFF;
    'h004018B4:rddata=8'h0F;
    'h004018B5:rddata=8'h0F;
    'h004018B6:rddata=8'h83;
    'h004018B7:rddata=8'h3D;
    'h004018B8:rddata=8'hFC;
    'h004018B9:rddata=8'h66;
    'h004018BA:rddata=8'h50;
    'h004018BB:rddata=8'h66;
    'h004018BC:rddata=8'h83;
    'h004018BD:rddata=8'hE8;
    'h004018BE:rddata=8'h02;
    'h004018BF:rddata=8'h66;
    'h004018C0:rddata=8'h0F;
    'h004018C1:rddata=8'hB6;
    'h004018C2:rddata=8'h5E;
    'h004018C3:rddata=8'h0D;
    'h004018C4:rddata=8'h8B;
    'h004018C5:rddata=8'hF3;
    'h004018C6:rddata=8'h66;
    'h004018C7:rddata=8'hF7;
    'h004018C8:rddata=8'hE3;
    'h004018C9:rddata=8'h66;
    'h004018CA:rddata=8'h03;
    'h004018CB:rddata=8'h46;
    'h004018CC:rddata=8'hFC;
    'h004018CD:rddata=8'hBB;
    'h004018CF:rddata=8'h82;
    'h004018D0:rddata=8'h8B;
    'h004018D1:rddata=8'hFB;
    'h004018D2:rddata=8'hB9;
    'h004018D3:rddata=8'h01;
    'h004018D5:rddata=8'hE8;
    'h004018D6:rddata=8'h28;
    'h004018D7:rddata=8'hFC;
    'h004018D8:rddata=8'h38;
    'h004018D9:rddata=8'h2D;
    'h004018DA:rddata=8'h74;
    'h004018DB:rddata=8'h1E;
    'h004018DC:rddata=8'hB1;
    'h004018DD:rddata=8'h0B;
    'h004018DE:rddata=8'h56;
    'h004018DF:rddata=8'hBE;
    'h004018E0:rddata=8'h6D;
    'h004018E1:rddata=8'h7D;
    'h004018E2:rddata=8'hF3;
    'h004018E3:rddata=8'hA6;
    'h004018E4:rddata=8'h5E;
    'h004018E5:rddata=8'h74;
    'h004018E6:rddata=8'h1B;
    'h004018E7:rddata=8'h03;
    'h004018E8:rddata=8'hF9;
    'h004018E9:rddata=8'h83;
    'h004018EA:rddata=8'hC7;
    'h004018EB:rddata=8'h15;
    'h004018EC:rddata=8'h3B;
    'h004018ED:rddata=8'hFB;
    'h004018EE:rddata=8'h72;
    'h004018EF:rddata=8'hE8;
    'h004018F0:rddata=8'h4E;
    'h004018F1:rddata=8'h75;
    'h004018F2:rddata=8'hDA;
    'h004018F3:rddata=8'h66;
    'h004018F4:rddata=8'h58;
    'h004018F5:rddata=8'hE8;
    'h004018F6:rddata=8'h65;
    'h004018F8:rddata=8'h72;
    'h004018F9:rddata=8'hBF;
    'h004018FA:rddata=8'h83;
    'h004018FB:rddata=8'hC4;
    'h004018FC:rddata=8'h04;
    'h004018FD:rddata=8'hE9;
    'h004018FE:rddata=8'hF6;
    'h004018FF:rddata=8'hFB;
    'h00401901:rddata=8'h20;
    'h00401902:rddata=8'h83;
    'h00401903:rddata=8'hC4;
    'h00401904:rddata=8'h04;
    'h00401905:rddata=8'h8B;
    'h00401906:rddata=8'h75;
    'h00401907:rddata=8'h09;
    'h00401908:rddata=8'h8B;
    'h00401909:rddata=8'h7D;
    'h0040190A:rddata=8'h0F;
    'h0040190B:rddata=8'h8B;
    'h0040190C:rddata=8'hC6;
    'h0040190D:rddata=8'h66;
    'h0040190E:rddata=8'hC1;
    'h0040190F:rddata=8'hE0;
    'h00401910:rddata=8'h10;
    'h00401911:rddata=8'h8B;
    'h00401912:rddata=8'hC7;
    'h00401913:rddata=8'h66;
    'h00401914:rddata=8'h83;
    'h00401915:rddata=8'hF8;
    'h00401916:rddata=8'h02;
    'h00401917:rddata=8'h0F;
    'h00401918:rddata=8'h82;
    'h00401919:rddata=8'hDB;
    'h0040191A:rddata=8'hFB;
    'h0040191B:rddata=8'h66;
    'h0040191C:rddata=8'h3D;
    'h0040191D:rddata=8'hF8;
    'h0040191E:rddata=8'hFF;
    'h0040191F:rddata=8'hFF;
    'h00401920:rddata=8'h0F;
    'h00401921:rddata=8'h0F;
    'h00401922:rddata=8'h83;
    'h00401923:rddata=8'hD1;
    'h00401924:rddata=8'hFB;
    'h00401925:rddata=8'h66;
    'h00401926:rddata=8'h50;
    'h00401927:rddata=8'h66;
    'h00401928:rddata=8'h83;
    'h00401929:rddata=8'hE8;
    'h0040192A:rddata=8'h02;
    'h0040192B:rddata=8'h66;
    'h0040192C:rddata=8'h0F;
    'h0040192D:rddata=8'hB6;
    'h0040192E:rddata=8'h4E;
    'h0040192F:rddata=8'h0D;
    'h00401930:rddata=8'h66;
    'h00401931:rddata=8'hF7;
    'h00401932:rddata=8'hE1;
    'h00401933:rddata=8'h66;
    'h00401934:rddata=8'h03;
    'h00401935:rddata=8'h46;
    'h00401936:rddata=8'hFC;
    'h00401937:rddata=8'hBB;
    'h0040193A:rddata=8'h06;
    'h0040193B:rddata=8'h8E;
    'h0040193C:rddata=8'h06;
    'h0040193E:rddata=8'h81;
    'h0040193F:rddata=8'hE8;
    'h00401940:rddata=8'hBE;
    'h00401941:rddata=8'hFB;
    'h00401942:rddata=8'h07;
    'h00401943:rddata=8'h66;
    'h00401944:rddata=8'h58;
    'h00401945:rddata=8'hC1;
    'h00401946:rddata=8'hEB;
    'h00401947:rddata=8'h04;
    'h00401948:rddata=8'h01;
    'h00401949:rddata=8'h1E;
    'h0040194B:rddata=8'h81;
    'h0040194C:rddata=8'hE8;
    'h0040194D:rddata=8'h0E;
    'h0040194F:rddata=8'h0F;
    'h00401950:rddata=8'h83;
    'h00401951:rddata=8'h02;
    'h00401953:rddata=8'h72;
    'h00401954:rddata=8'hD0;
    'h00401955:rddata=8'h8A;
    'h00401956:rddata=8'h56;
    'h00401957:rddata=8'h40;
    'h00401958:rddata=8'hEA;
    'h0040195C:rddata=8'h20;
    'h0040195D:rddata=8'h66;
    'h0040195E:rddata=8'hC1;
    'h0040195F:rddata=8'hE0;
    'h00401960:rddata=8'h02;
    'h00401961:rddata=8'hE8;
    'h00401962:rddata=8'h11;
    'h00401964:rddata=8'h26;
    'h00401965:rddata=8'h66;
    'h00401966:rddata=8'h8B;
    'h00401967:rddata=8'h01;
    'h00401968:rddata=8'h66;
    'h00401969:rddata=8'h25;
    'h0040196A:rddata=8'hFF;
    'h0040196B:rddata=8'hFF;
    'h0040196C:rddata=8'hFF;
    'h0040196D:rddata=8'h0F;
    'h0040196E:rddata=8'h66;
    'h0040196F:rddata=8'h3D;
    'h00401970:rddata=8'hF8;
    'h00401971:rddata=8'hFF;
    'h00401972:rddata=8'hFF;
    'h00401973:rddata=8'h0F;
    'h00401974:rddata=8'hC3;
    'h00401975:rddata=8'hBF;
    'h00401977:rddata=8'h7E;
    'h00401978:rddata=8'h66;
    'h00401979:rddata=8'h0F;
    'h0040197A:rddata=8'hB7;
    'h0040197B:rddata=8'h4E;
    'h0040197C:rddata=8'h0B;
    'h0040197D:rddata=8'h66;
    'h0040197E:rddata=8'h33;
    'h0040197F:rddata=8'hD2;
    'h00401980:rddata=8'h66;
    'h00401981:rddata=8'hF7;
    'h00401982:rddata=8'hF1;
    'h00401983:rddata=8'h66;
    'h00401984:rddata=8'h3B;
    'h00401985:rddata=8'h46;
    'h00401986:rddata=8'hF4;
    'h00401987:rddata=8'h74;
    'h00401988:rddata=8'h3A;
    'h00401989:rddata=8'h66;
    'h0040198A:rddata=8'h89;
    'h0040198B:rddata=8'h46;
    'h0040198C:rddata=8'hF4;
    'h0040198D:rddata=8'h66;
    'h0040198E:rddata=8'h03;
    'h0040198F:rddata=8'h46;
    'h00401990:rddata=8'h1C;
    'h00401991:rddata=8'h66;
    'h00401992:rddata=8'h0F;
    'h00401993:rddata=8'hB7;
    'h00401994:rddata=8'h4E;
    'h00401995:rddata=8'h0E;
    'h00401996:rddata=8'h66;
    'h00401997:rddata=8'h03;
    'h00401998:rddata=8'hC1;
    'h00401999:rddata=8'h66;
    'h0040199A:rddata=8'h0F;
    'h0040199B:rddata=8'hB7;
    'h0040199C:rddata=8'h5E;
    'h0040199D:rddata=8'h28;
    'h0040199E:rddata=8'h83;
    'h0040199F:rddata=8'hE3;
    'h004019A0:rddata=8'h0F;
    'h004019A1:rddata=8'h74;
    'h004019A2:rddata=8'h16;
    'h004019A3:rddata=8'h3A;
    'h004019A4:rddata=8'h5E;
    'h004019A5:rddata=8'h10;
    'h004019A6:rddata=8'h0F;
    'h004019A7:rddata=8'h83;
    'h004019A8:rddata=8'h4C;
    'h004019A9:rddata=8'hFB;
    'h004019AA:rddata=8'h52;
    'h004019AB:rddata=8'h66;
    'h004019AC:rddata=8'h8B;
    'h004019AD:rddata=8'hC8;
    'h004019AE:rddata=8'h66;
    'h004019AF:rddata=8'h8B;
    'h004019B0:rddata=8'h46;
    'h004019B1:rddata=8'h24;
    'h004019B2:rddata=8'h66;
    'h004019B3:rddata=8'hF7;
    'h004019B4:rddata=8'hE3;
    'h004019B5:rddata=8'h66;
    'h004019B6:rddata=8'h03;
    'h004019B7:rddata=8'hC1;
    'h004019B8:rddata=8'h5A;
    'h004019B9:rddata=8'h52;
    'h004019BA:rddata=8'h8B;
    'h004019BB:rddata=8'hDF;
    'h004019BC:rddata=8'hB9;
    'h004019BD:rddata=8'h01;
    'h004019BF:rddata=8'hE8;
    'h004019C0:rddata=8'h3E;
    'h004019C1:rddata=8'hFB;
    'h004019C2:rddata=8'h5A;
    'h004019C3:rddata=8'h8B;
    'h004019C4:rddata=8'hDA;
    'h004019C5:rddata=8'hC3;
    'h004019FE:rddata=8'h55;
    'h004019FF:rddata=8'hAA;
    'h00632800:rddata=8'hF8;
    'h00632801:rddata=8'hFF;
    'h00632802:rddata=8'hFF;
    'h00632803:rddata=8'h0F;
    'h00632804:rddata=8'hFF;
    'h00632805:rddata=8'hFF;
    'h00632806:rddata=8'hFF;
    'h00632807:rddata=8'hFF;
    'h00632808:rddata=8'hFF;
    'h00632809:rddata=8'hFF;
    'h0063280A:rddata=8'hFF;
    'h0063280B:rddata=8'h0F;
    'h0063280C:rddata=8'hFF;
    'h0063280D:rddata=8'hFF;
    'h0063280E:rddata=8'hFF;
    'h0063280F:rddata=8'h0F;
    'h00632810:rddata=8'hFF;
    'h00632811:rddata=8'hFF;
    'h00632812:rddata=8'hFF;
    'h00632813:rddata=8'h0F;
    'h00632814:rddata=8'hFF;
    'h00632815:rddata=8'hFF;
    'h00632816:rddata=8'hFF;
    'h00632817:rddata=8'h0F;
    'h00632818:rddata=8'hFF;
    'h00632819:rddata=8'hFF;
    'h0063281A:rddata=8'hFF;
    'h0063281B:rddata=8'h0F;
    'h00719400:rddata=8'hF8;
    'h00719401:rddata=8'hFF;
    'h00719402:rddata=8'hFF;
    'h00719403:rddata=8'h0F;
    'h00719404:rddata=8'hFF;
    'h00719405:rddata=8'hFF;
    'h00719406:rddata=8'hFF;
    'h00719407:rddata=8'hFF;
    'h00719408:rddata=8'hFF;
    'h00719409:rddata=8'hFF;
    'h0071940A:rddata=8'hFF;
    'h0071940B:rddata=8'h0F;
    'h0071940C:rddata=8'hFF;
    'h0071940D:rddata=8'hFF;
    'h0071940E:rddata=8'hFF;
    'h0071940F:rddata=8'h0F;
    'h00719410:rddata=8'hFF;
    'h00719411:rddata=8'hFF;
    'h00719412:rddata=8'hFF;
    'h00719413:rddata=8'h0F;
    'h00719414:rddata=8'hFF;
    'h00719415:rddata=8'hFF;
    'h00719416:rddata=8'hFF;
    'h00719417:rddata=8'h0F;
    'h00719418:rddata=8'hFF;
    'h00719419:rddata=8'hFF;
    'h0071941A:rddata=8'hFF;
    'h0071941B:rddata=8'h0F;
    'h00800000:rddata=8'h42;
    'h00800001:rddata=8'h20;
    'h00800003:rddata=8'h49;
    'h00800005:rddata=8'h6E;
    'h00800007:rddata=8'h66;
    'h00800009:rddata=8'h6F;
    'h0080000B:rddata=8'h0F;
    'h0080000D:rddata=8'h72;
    'h0080000E:rddata=8'h72;
    'h00800010:rddata=8'h6D;
    'h00800012:rddata=8'h61;
    'h00800014:rddata=8'h74;
    'h00800016:rddata=8'h69;
    'h00800018:rddata=8'h6F;
    'h0080001C:rddata=8'h6E;
    'h00800020:rddata=8'h01;
    'h00800021:rddata=8'h53;
    'h00800023:rddata=8'h79;
    'h00800025:rddata=8'h73;
    'h00800027:rddata=8'h74;
    'h00800029:rddata=8'h65;
    'h0080002B:rddata=8'h0F;
    'h0080002D:rddata=8'h72;
    'h0080002E:rddata=8'h6D;
    'h00800030:rddata=8'h20;
    'h00800032:rddata=8'h56;
    'h00800034:rddata=8'h6F;
    'h00800036:rddata=8'h6C;
    'h00800038:rddata=8'h75;
    'h0080003C:rddata=8'h6D;
    'h0080003E:rddata=8'h65;
    'h00800040:rddata=8'h53;
    'h00800041:rddata=8'h59;
    'h00800042:rddata=8'h53;
    'h00800043:rddata=8'h54;
    'h00800044:rddata=8'h45;
    'h00800045:rddata=8'h4D;
    'h00800046:rddata=8'h7E;
    'h00800047:rddata=8'h31;
    'h00800048:rddata=8'h20;
    'h00800049:rddata=8'h20;
    'h0080004A:rddata=8'h20;
    'h0080004B:rddata=8'h16;
    'h0080004D:rddata=8'h69;
    'h0080004E:rddata=8'h7C;
    'h0080004F:rddata=8'h0A;
    'h00800050:rddata=8'hE4;
    'h00800051:rddata=8'h4E;
    'h00800052:rddata=8'hE4;
    'h00800053:rddata=8'h4E;
    'h00800056:rddata=8'h7D;
    'h00800057:rddata=8'h0A;
    'h00800058:rddata=8'hE4;
    'h00800059:rddata=8'h4E;
    'h0080005A:rddata=8'h03;
    'h00800060:rddata=8'hE5;
    'h00800061:rddata=8'hB0;
    'h00800062:rddata=8'h65;
    'h00800063:rddata=8'hFA;
    'h00800064:rddata=8'h5E;
    'h00800065:rddata=8'h87;
    'h00800066:rddata=8'h65;
    'h00800067:rddata=8'h2C;
    'h00800068:rddata=8'h67;
    'h00800069:rddata=8'h87;
    'h0080006A:rddata=8'h65;
    'h0080006B:rddata=8'h0F;
    'h0080006D:rddata=8'hD2;
    'h0080006E:rddata=8'h63;
    'h0080006F:rddata=8'h68;
    'h00800070:rddata=8'h2E;
    'h00800072:rddata=8'h74;
    'h00800074:rddata=8'h78;
    'h00800076:rddata=8'h74;
    'h0080007C:rddata=8'hFF;
    'h0080007D:rddata=8'hFF;
    'h0080007E:rddata=8'hFF;
    'h0080007F:rddata=8'hFF;
    'h00800080:rddata=8'hE5;
    'h00800081:rddata=8'hC2;
    'h00800082:rddata=8'hBD;
    'h00800083:rddata=8'hA8;
    'h00800084:rddata=8'hCE;
    'h00800085:rddata=8'hC4;
    'h00800086:rddata=8'h7E;
    'h00800087:rddata=8'h31;
    'h00800088:rddata=8'h54;
    'h00800089:rddata=8'h58;
    'h0080008A:rddata=8'h54;
    'h0080008B:rddata=8'h20;
    'h0080008D:rddata=8'h5C;
    'h0080008E:rddata=8'hD4;
    'h0080008F:rddata=8'h0A;
    'h00800090:rddata=8'hE4;
    'h00800091:rddata=8'h4E;
    'h00800092:rddata=8'hE4;
    'h00800093:rddata=8'h4E;
    'h00800096:rddata=8'hD5;
    'h00800097:rddata=8'h0A;
    'h00800098:rddata=8'hE4;
    'h00800099:rddata=8'h4E;
    'h008000A0:rddata=8'h42;
    'h008000A1:rddata=8'h53;
    'h008000A3:rddata=8'h44;
    'h008000A5:rddata=8'h63;
    'h008000A7:rddata=8'h61;
    'h008000A9:rddata=8'h72;
    'h008000AB:rddata=8'h0F;
    'h008000AD:rddata=8'h9F;
    'h008000AE:rddata=8'h64;
    'h008000B0:rddata=8'h2E;
    'h008000B2:rddata=8'h74;
    'h008000B4:rddata=8'h78;
    'h008000B6:rddata=8'h74;
    'h008000BC:rddata=8'hFF;
    'h008000BD:rddata=8'hFF;
    'h008000BE:rddata=8'hFF;
    'h008000BF:rddata=8'hFF;
    'h008000C0:rddata=8'h01;
    'h008000C1:rddata=8'h46;
    'h008000C3:rddata=8'h69;
    'h008000C5:rddata=8'h6C;
    'h008000C7:rddata=8'h65;
    'h008000C9:rddata=8'h2D;
    'h008000CB:rddata=8'h0F;
    'h008000CD:rddata=8'h9F;
    'h008000CE:rddata=8'h69;
    'h008000D0:rddata=8'h6E;
    'h008000D2:rddata=8'h2D;
    'h008000D4:rddata=8'h66;
    'h008000D6:rddata=8'h61;
    'h008000D8:rddata=8'h6B;
    'h008000DC:rddata=8'h65;
    'h008000DE:rddata=8'h2D;
    'h008000E0:rddata=8'h46;
    'h008000E1:rddata=8'h49;
    'h008000E2:rddata=8'h4C;
    'h008000E3:rddata=8'h45;
    'h008000E4:rddata=8'h2D;
    'h008000E5:rddata=8'h49;
    'h008000E6:rddata=8'h7E;
    'h008000E7:rddata=8'h31;
    'h008000E8:rddata=8'h54;
    'h008000E9:rddata=8'h58;
    'h008000EA:rddata=8'h54;
    'h008000EB:rddata=8'h20;
    'h008000ED:rddata=8'h5C;
    'h008000EE:rddata=8'hD4;
    'h008000EF:rddata=8'h0A;
    'h008000F0:rddata=8'hE4;
    'h008000F1:rddata=8'h4E;
    'h008000F2:rddata=8'hE4;
    'h008000F3:rddata=8'h4E;
    'h008000F6:rddata=8'hF0;
    'h008000F7:rddata=8'h0A;
    'h008000F8:rddata=8'hE4;
    'h008000F9:rddata=8'h4E;
    'h008000FA:rddata=8'h06;
    'h008000FC:rddata=8'h12;
    'h00808000:rddata=8'h2E;
    'h00808001:rddata=8'h20;
    'h00808002:rddata=8'h20;
    'h00808003:rddata=8'h20;
    'h00808004:rddata=8'h20;
    'h00808005:rddata=8'h20;
    'h00808006:rddata=8'h20;
    'h00808007:rddata=8'h20;
    'h00808008:rddata=8'h20;
    'h00808009:rddata=8'h20;
    'h0080800A:rddata=8'h20;
    'h0080800B:rddata=8'h10;
    'h0080800D:rddata=8'h69;
    'h0080800E:rddata=8'h7C;
    'h0080800F:rddata=8'h0A;
    'h00808010:rddata=8'hE4;
    'h00808011:rddata=8'h4E;
    'h00808012:rddata=8'hE4;
    'h00808013:rddata=8'h4E;
    'h00808016:rddata=8'h7D;
    'h00808017:rddata=8'h0A;
    'h00808018:rddata=8'hE4;
    'h00808019:rddata=8'h4E;
    'h0080801A:rddata=8'h03;
    'h00808020:rddata=8'h2E;
    'h00808021:rddata=8'h2E;
    'h00808022:rddata=8'h20;
    'h00808023:rddata=8'h20;
    'h00808024:rddata=8'h20;
    'h00808025:rddata=8'h20;
    'h00808026:rddata=8'h20;
    'h00808027:rddata=8'h20;
    'h00808028:rddata=8'h20;
    'h00808029:rddata=8'h20;
    'h0080802A:rddata=8'h20;
    'h0080802B:rddata=8'h10;
    'h0080802D:rddata=8'h69;
    'h0080802E:rddata=8'h7C;
    'h0080802F:rddata=8'h0A;
    'h00808030:rddata=8'hE4;
    'h00808031:rddata=8'h4E;
    'h00808032:rddata=8'hE4;
    'h00808033:rddata=8'h4E;
    'h00808036:rddata=8'h7D;
    'h00808037:rddata=8'h0A;
    'h00808038:rddata=8'hE4;
    'h00808039:rddata=8'h4E;
    'h00808040:rddata=8'h42;
    'h00808041:rddata=8'h74;
    'h00808045:rddata=8'hFF;
    'h00808046:rddata=8'hFF;
    'h00808047:rddata=8'hFF;
    'h00808048:rddata=8'hFF;
    'h00808049:rddata=8'hFF;
    'h0080804A:rddata=8'hFF;
    'h0080804B:rddata=8'h0F;
    'h0080804D:rddata=8'hCE;
    'h0080804E:rddata=8'hFF;
    'h0080804F:rddata=8'hFF;
    'h00808050:rddata=8'hFF;
    'h00808051:rddata=8'hFF;
    'h00808052:rddata=8'hFF;
    'h00808053:rddata=8'hFF;
    'h00808054:rddata=8'hFF;
    'h00808055:rddata=8'hFF;
    'h00808056:rddata=8'hFF;
    'h00808057:rddata=8'hFF;
    'h00808058:rddata=8'hFF;
    'h00808059:rddata=8'hFF;
    'h0080805C:rddata=8'hFF;
    'h0080805D:rddata=8'hFF;
    'h0080805E:rddata=8'hFF;
    'h0080805F:rddata=8'hFF;
    'h00808060:rddata=8'h01;
    'h00808061:rddata=8'h57;
    'h00808063:rddata=8'h50;
    'h00808065:rddata=8'h53;
    'h00808067:rddata=8'h65;
    'h00808069:rddata=8'h74;
    'h0080806B:rddata=8'h0F;
    'h0080806D:rddata=8'hCE;
    'h0080806E:rddata=8'h74;
    'h00808070:rddata=8'h69;
    'h00808072:rddata=8'h6E;
    'h00808074:rddata=8'h67;
    'h00808076:rddata=8'h73;
    'h00808078:rddata=8'h2E;
    'h0080807C:rddata=8'h64;
    'h0080807E:rddata=8'h61;
    'h00808080:rddata=8'h57;
    'h00808081:rddata=8'h50;
    'h00808082:rddata=8'h53;
    'h00808083:rddata=8'h45;
    'h00808084:rddata=8'h54;
    'h00808085:rddata=8'h54;
    'h00808086:rddata=8'h7E;
    'h00808087:rddata=8'h31;
    'h00808088:rddata=8'h44;
    'h00808089:rddata=8'h41;
    'h0080808A:rddata=8'h54;
    'h0080808B:rddata=8'h20;
    'h0080808D:rddata=8'h73;
    'h0080808E:rddata=8'h7C;
    'h0080808F:rddata=8'h0A;
    'h00808090:rddata=8'hE4;
    'h00808091:rddata=8'h4E;
    'h00808092:rddata=8'hE4;
    'h00808093:rddata=8'h4E;
    'h00808096:rddata=8'h7D;
    'h00808097:rddata=8'h0A;
    'h00808098:rddata=8'hE4;
    'h00808099:rddata=8'h4E;
    'h0080809A:rddata=8'h04;
    'h0080809C:rddata=8'h0C;
    'h008080A0:rddata=8'h42;
    'h008080A1:rddata=8'h47;
    'h008080A3:rddata=8'h75;
    'h008080A5:rddata=8'h69;
    'h008080A7:rddata=8'h64;
    'h008080AB:rddata=8'h0F;
    'h008080AD:rddata=8'hFF;
    'h008080AE:rddata=8'hFF;
    'h008080AF:rddata=8'hFF;
    'h008080B0:rddata=8'hFF;
    'h008080B1:rddata=8'hFF;
    'h008080B2:rddata=8'hFF;
    'h008080B3:rddata=8'hFF;
    'h008080B4:rddata=8'hFF;
    'h008080B5:rddata=8'hFF;
    'h008080B6:rddata=8'hFF;
    'h008080B7:rddata=8'hFF;
    'h008080B8:rddata=8'hFF;
    'h008080B9:rddata=8'hFF;
    'h008080BC:rddata=8'hFF;
    'h008080BD:rddata=8'hFF;
    'h008080BE:rddata=8'hFF;
    'h008080BF:rddata=8'hFF;
    'h008080C0:rddata=8'h01;
    'h008080C1:rddata=8'h49;
    'h008080C3:rddata=8'h6E;
    'h008080C5:rddata=8'h64;
    'h008080C7:rddata=8'h65;
    'h008080C9:rddata=8'h78;
    'h008080CB:rddata=8'h0F;
    'h008080CD:rddata=8'hFF;
    'h008080CE:rddata=8'h65;
    'h008080D0:rddata=8'h72;
    'h008080D2:rddata=8'h56;
    'h008080D4:rddata=8'h6F;
    'h008080D6:rddata=8'h6C;
    'h008080D8:rddata=8'h75;
    'h008080DC:rddata=8'h6D;
    'h008080DE:rddata=8'h65;
    'h008080E0:rddata=8'h49;
    'h008080E1:rddata=8'h4E;
    'h008080E2:rddata=8'h44;
    'h008080E3:rddata=8'h45;
    'h008080E4:rddata=8'h58;
    'h008080E5:rddata=8'h45;
    'h008080E6:rddata=8'h7E;
    'h008080E7:rddata=8'h31;
    'h008080E8:rddata=8'h20;
    'h008080E9:rddata=8'h20;
    'h008080EA:rddata=8'h20;
    'h008080EB:rddata=8'h20;
    'h008080ED:rddata=8'h31;
    'h008080EE:rddata=8'h80;
    'h008080EF:rddata=8'h0A;
    'h008080F0:rddata=8'hE4;
    'h008080F1:rddata=8'h4E;
    'h008080F2:rddata=8'hE4;
    'h008080F3:rddata=8'h4E;
    'h008080F6:rddata=8'h81;
    'h008080F7:rddata=8'h0A;
    'h008080F8:rddata=8'hE4;
    'h008080F9:rddata=8'h4E;
    'h008080FA:rddata=8'h05;
    'h008080FC:rddata=8'h4C;
    'h00818000:rddata=8'h7B;
    'h00818002:rddata=8'h30;
    'h00818004:rddata=8'h41;
    'h00818006:rddata=8'h30;
    'h00818008:rddata=8'h39;
    'h0081800A:rddata=8'h42;
    'h0081800C:rddata=8'h35;
    'h0081800E:rddata=8'h39;
    'h00818010:rddata=8'h34;
    'h00818012:rddata=8'h2D;
    'h00818014:rddata=8'h33;
    'h00818016:rddata=8'h34;
    'h00818018:rddata=8'h45;
    'h0081801A:rddata=8'h35;
    'h0081801C:rddata=8'h2D;
    'h0081801E:rddata=8'h34;
    'h00818020:rddata=8'h33;
    'h00818022:rddata=8'h41;
    'h00818024:rddata=8'h43;
    'h00818026:rddata=8'h2D;
    'h00818028:rddata=8'h38;
    'h0081802A:rddata=8'h30;
    'h0081802C:rddata=8'h35;
    'h0081802E:rddata=8'h44;
    'h00818030:rddata=8'h2D;
    'h00818032:rddata=8'h43;
    'h00818034:rddata=8'h32;
    'h00818036:rddata=8'h30;
    'h00818038:rddata=8'h43;
    'h0081803A:rddata=8'h30;
    'h0081803C:rddata=8'h39;
    'h0081803E:rddata=8'h36;
    'h00818040:rddata=8'h36;
    'h00818042:rddata=8'h37;
    'h00818044:rddata=8'h31;
    'h00818046:rddata=8'h41;
    'h00818048:rddata=8'h31;
    'h0081804A:rddata=8'h7D;
    'h00810000:rddata=8'h0C;
    'h00810004:rddata=8'hB7;
    'h00810005:rddata=8'hF3;
    'h00810006:rddata=8'hA4;
    'h00810007:rddata=8'h26;
    'h00810008:rddata=8'h3D;
    'h00810009:rddata=8'hE2;
    'h0081000A:rddata=8'h84;
    'h0081000B:rddata=8'h39;
    'h00820000:rddata=8'h49;
    'h00820001:rddata=8'h27;
    'h00820002:rddata=8'h6D;
    'h00820003:rddata=8'h20;
    'h00820004:rddata=8'h61;
    'h00820005:rddata=8'h20;
    'h00820006:rddata=8'h66;
    'h00820007:rddata=8'h61;
    'h00820008:rddata=8'h6B;
    'h00820009:rddata=8'h65;
    'h0082000A:rddata=8'h20;
    'h0082000B:rddata=8'h73;
    'h0082000C:rddata=8'h64;
    'h0082000D:rddata=8'h63;
    'h0082000E:rddata=8'h61;
    'h0082000F:rddata=8'h72;
    'h00820010:rddata=8'h64;
    'h00820011:rddata=8'h21;
    default   :rddata=8'h00;
    endcase

endmodule
